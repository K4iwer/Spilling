module roberto_uc (
    input wire clock,
    input wire reset,
    input wire pronto_medida1,
    input wire pronto_medida2,
    input wire pronto_medida3,
    
)





endmodule